//countervar_v1_tb.sv by Vincent Gosselin,2020.
//testbench in SystemVerilog for variable counter up / down 

// input free_time;

// free_time = 1;

// while(free_time) begin
	// $display ("continue to pwn");
// end